 //Top Level Module for Traffic Lights Project
module traffic_lights(
		//Input Wires
		input wire clk, //Clock signal, from Crystal Oscillator on board 
		input wire reset, //Reset signal, triggered by user by pressing physical button
		input wire pedestrian, //Signal to simulate pedestrian crossing road, physical button
		//Output Wires
		output wire Red, //If HIGH (1), the red light will be lit 
		output wire Amber, //If HIGH (1), the amber light will be lit
		output wire Green, //If HIGH (1), the green light will be lit 
		output wire Flag //If HIGH (1), an LED will be lit to show pedestrian state				
    );
	 
	localparam scale_to_second = 25000000; //Parameter to scale Crystal Oscillator Frequency 
										  //to 1 second period
	wire second_clk; //Wire to carry the 1Hz clock signal between modules, as generated by the 
					//scaled frequency
	wire[3:0] counter; //Wire to carry the value of the counter between modules, 4bits wide
	wire[1:0] curr_colour;	//Wire to carry the value of the current light colour between modules, 
							//2bits wide
	wire red_wire, amber_wire, green_wire; //Wires to carry signal for light to be lit, 
										   //give output to module
	wire ped_wire; //Wire to carry signal for pedestrian indicator LED
	
	//Instantiate the clock module to provide 1Hz clock signal
	clock clk_second(.CCLK(clk), .clkscale(scale_to_second), .clk(second_clk));
	
	//Instantiate the counter to keep track of how long the current colour has been lit (curr_colour)
	light_timer timing(.clk(second_clk), .reset(reset), .curr_code(curr_colour), .timer_reg(counter));
	
	//Instantiate the control module to decide which state we are in and which light should be lit
	lights_control controller(.clk(second_clk), .ped_flag_in(ped_wire), .reset(reset), 
			.pedestrian(pedestrian), .count(counter), .state_reg(curr_colour), .ped_flag_out(ped_wire));
	
	//Instantiate the multiplexer module to enable assigning of light to be lit, based on output 
	//of the control module
	multiplexer choice(.colour_code(curr_colour), .red_reg(red_wire), 
						.amber_reg(amber_wire), .green_reg(green_wire));
	
	//Assignments of lights to be lit
	assign Red = red_wire;
	assign Amber = amber_wire;
	assign Green = green_wire;
	assign Flag = ped_wire;
	
endmodule